`define SCREEN_WIDTH 176
`define SCREEN_HEIGHT 144

module IMAGE_PROCESSOR (

);


//=======================================================
//  PARAMETER declarations
//=======================================================


//=======================================================
//  PORT declarations
//=======================================================


//=======================================================
//  PROCESSING
//=======================================================


endmodule